module uart_top #() ();


    // UART TXR

    // UART RXR

    // UART FIFO

    // UART BUAD_GENERATOR
    
endmodule : uart_top